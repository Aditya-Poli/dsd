/* AND Gate Gate Level Modelling
   This file conatains AND Gate module
   using Gate Level Modelling
*/

module AND_GLM(output Y, input A, B);
    and(Y, A, B);
endmodule